module FullAdder_4Bit(i_1, i_2, i_c, o_s, o_c);

    input [4:0]i_1, [4:0]i_2, [4:0]i_c;
    output [4:0]o_s, o_c;
    wire [3:0]o_cw;

    

endmodule